module char_rom (
input logic [5:0] rom_address, // 16 addresses in total
output logic [63:0] rom_data); // 64bits/address

always_comb

begin
case (rom_address)
6'b000000 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000001 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000010 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000011 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000100 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000101 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000110 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b000111 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b001000 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100101 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100110 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100111 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101000 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101001 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101010 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101011 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b001001 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b001010 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b001011 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b001100 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b001101 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b001110 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b001111 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b010000 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b010001 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b010010 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b010011 : rom_data = 64'b1111111111111111111111100000000000000000111111111111111111111111;
6'b010100 : rom_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
6'b010101 : rom_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
6'b010110 : rom_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
6'b010111 : rom_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
6'b011000 : rom_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
6'b011001 : rom_data = 64'b1111111111111111111111100000000000000001111111111111111111111111;
6'b011010 : rom_data = 64'b1111111111111111111111100000000000000001111111111111111111111111;
6'b011011 : rom_data = 64'b1111111111111111111111100000000000000001111111111111111111111111;
6'b011100 : rom_data = 64'b1111111111111111111111100000000000000001111111111111111111111111;
6'b011101 : rom_data = 64'b1111111111111111111111100000000000000001111111111111111111111111;
6'b011110 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b011111 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100000 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100001 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100010 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100011 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b100100 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101100 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101101 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101110 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'b101111 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
default	 : rom_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
endcase;

end

endmodule
